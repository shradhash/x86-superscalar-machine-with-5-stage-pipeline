package CACHE;

typedef enum {IDLE,
              READ,
              WRITE,
              FLUSH} req_type;

endpackage

